* netlist generated with vector fitting poles and residues

.subckt total_network node_1 node_2 node_3 node_4 node_ref
X_11 node_1 node_ref yp11
X_12 node_1 node_2 yp12
X_13 node_1 node_3 yp13
X_14 node_1 node_4 yp14
X_22 node_2 node_ref yp22
X_23 node_2 node_3 yp23
X_24 node_2 node_4 yp24
X_33 node_3 node_ref yp33
X_34 node_3 node_4 yp34
X_44 node_4 node_ref yp44
.ends


* Y'11
.subckt yp11 node_1 node_ref
* Branch 0
Rabr0 node_1 netRa0 1019.5086409595948
Lbr0 netRa0 netL0 1.7666142776744992e-07
Rbbr0 netL0 node_ref -197.5274565119536
Cbr0 netL0 node_ref 9.254922024746562e-13

* Branch 1
Rabr1 node_1 netRa1 -1461.7244879191398
Lbr1 netRa1 netL1 1.3330432121141119e-06
Rbbr1 netL1 node_ref -38046.92323675643
Cbr1 netL1 node_ref 1.8283307991714893e-14

* Branch 2
Rabr2 node_1 netRa2 24.235729720999508
Lbr2 netRa2 netL2 1.7825337242182876e-07
Rbbr2 netL2 node_ref -145808.3659864874
Cbr2 netL2 node_ref 1.4212847239721875e-13

* Branch 3
Rabr3 node_1 netRa3 41.2288276456704
Lbr3 netRa3 netL3 3.847071333987913e-07
Rbbr3 netL3 node_ref -21679.458849925693
Cbr3 netL3 node_ref 6.58659603468876e-14

* Branch 4
Rabr4 node_1 netRa4 -133.86328777920897
Lbr4 netRa4 netL4 2.5167302762380917e-07
Rbbr4 netL4 node_ref -3204.389551883395
Cbr4 netL4 node_ref 9.438874619745873e-14

* Branch 5
Rabr5 node_1 netRa5 -67118.42820570062
Lbr5 netRa5 netL5 3.285633153655026e-06
Rbbr5 netL5 node_ref -80621.06072223542
Cbr5 netL5 node_ref 4.362046050891356e-16

* Branch 6
Rabr6 node_1 netRa6 -12979.362978227513
Lbr6 netRa6 netL6 -2.984033700407258e-06
Rbbr6 netL6 node_ref -159853.1217332292
Cbr6 netL6 node_ref -1.9523301332220975e-15

* Branch 7
Rabr7 node_1 netRa7 8.320636551521098
Lbr7 netRa7 netL7 9.1288132070139e-08
Rbbr7 netL7 node_ref -34827.862277786444
Cbr7 netL7 node_ref 6.936967125319643e-14

* Branch 8
Rabr8 node_1 netRa8 24.716249057676055
Lbr8 netRa8 netL8 9.244064259689205e-08
Rbbr8 netL8 node_ref -4760.900255553137
Cbr8 netL8 node_ref 6.801646572955332e-14

* Branch 9
Rabr9 node_1 netRa9 683.3476830865044
Lbr9 netRa9 netL9 2.1950343237527242e-07
Rbbr9 netL9 node_ref 35034.86592871867
Cbr9 netL9 node_ref 1.2577346055400513e-14

* Branch 10
Rabr10 node_1 netRa10 -26.37796584651283
Lbr10 netRa10 netL10 5.974206365372397e-08
Rbbr10 netL10 node_ref -12566.746423558829
Cbr10 netL10 node_ref 4.6990039881431255e-14

* Branch 11
Rabr11 node_1 netRa11 -6100.774347545953
Lbr11 netRa11 netL11 -3.0778609219741427e-06
Rbbr11 netL11 node_ref 445842.6194710535
Cbr11 netL11 node_ref -5.356290379383056e-16

* Branch 12
Rabr12 node_1 netRa12 7670.559240469734
Lbr12 netRa12 netL12 9.988239779919354e-07
Rbbr12 netL12 node_ref 101931.55549203673
Cbr12 netL12 node_ref 1.4689394985549136e-15

* Branch 13
Rabr13 node_1 netRa13 -0.708841812375048
Lbr13 netRa13 netL13 3.9971163233651375e-08
Rbbr13 netL13 node_ref -15683.155190034424
Cbr13 netL13 node_ref 3.959783994475154e-14

* Branch 14
Rabr14 node_1 netRa14 3718.170231946571
Lbr14 netRa14 netL14 1.5527271011934648e-06
Rbbr14 netL14 node_ref 1543738.2984921318
Cbr14 netL14 node_ref 6.50169452562026e-16

* Branch 15
Rabr15 node_1 netRa15 -13.45156138419204
Lbr15 netRa15 netL15 3.394569179005267e-08
Rbbr15 netL15 node_ref -9853.489596117963
Cbr15 netL15 node_ref 2.9752975896587675e-14

* Branch 16
Rabr16 node_1 netRa16 -7.454793789419227
Lbr16 netRa16 netL16 9.624367778395192e-08
Rbbr16 netL16 node_ref -88962.47759269028
Cbr16 netL16 node_ref 7.312273775091523e-15

* Branch 17
Rabr17 node_1 netRa17 -250.24925291031326
Lbr17 netRa17 netL17 5.45170374213417e-08
Rbbr17 netL17 node_ref -9663.164902857188
Cbr17 netL17 node_ref 1.2468167730666732e-14

* Branch 18
Rabr18 node_1 netRa18 371.3040243462196
Lbr18 netRa18 netL18 1.2332205636415833e-08
Rbbr18 netL18 node_ref -516.6525134541523
Cbr18 netL18 node_ref 9.085708575877874e-14

* Branch 19
Rabr19 node_1 netRa19 -42.94757816236134
Lbr19 netRa19 netL19 7.186054054745924e-08
Rbbr19 netL19 node_ref -46666.4392101813
Cbr19 netL19 node_ref 7.187448290445781e-15

* Branch 20
Rabr20 node_1 netRa20 -2696.265596725878
Lbr20 netRa20 netL20 5.4148246381165245e-08
Rbbr20 netL20 node_ref -4614.755730212657
Cbr20 netL20 node_ref 3.724736640252133e-15

* Branch 21
Rabr21 node_1 netRa21 -373.5320034435647
Lbr21 netRa21 netL21 6.883274388317828e-08
Rbbr21 netL21 node_ref -20725.92389105796
Cbr21 netL21 node_ref 5.630037235937145e-15

* Branch 22
Rabr22 node_1 netRa22 126.33150651278649
Lbr22 netRa22 netL22 1.630396324756196e-08
Rbbr22 netL22 node_ref -7646.485123513112
Cbr22 netL22 node_ref 2.40676311164974e-14

* Branch 23
Rabr23 node_1 netRa23 87796.87367687559
Lbr23 netRa23 netL23 -6.035397745466925e-07
Rbbr23 netL23 node_ref 100504.98582246566
Cbr23 netL23 node_ref -6.561077863170135e-17

* Branch 24
Rabr24 node_1 netRa24 -77.3270105113985
Lbr24 netRa24 netL24 3.283496699416413e-08
Rbbr24 netL24 node_ref -20687.674519268905
Cbr24 netL24 node_ref 9.479905475564742e-15

.ends


* Y'12
.subckt yp12 node_1 node_2
* Branch 0
Rabr0 node_1 netRa0 -1860.8354455794627
Lbr0 netRa0 netL0 -2.829290628959974e-07
Rbbr0 netL0 node_2 425.1417295131353
Cbr0 netL0 node_2 -5.043117717297719e-13

* Branch 1
Rabr1 node_1 netRa1 -37.65479302274327
Lbr1 netRa1 netL1 -3.2433015793407737e-07
Rbbr1 netL1 node_2 56851.945071883565
Cbr1 netL1 node_2 -7.820118685330792e-14

* Branch 2
Rabr2 node_1 netRa2 -319.2672358827794
Lbr2 netRa2 netL2 -1.1484361081007304e-06
Rbbr2 netL2 node_2 -483740.9768089124
Cbr2 netL2 node_2 -2.204210650111845e-14

* Branch 3
Rabr3 node_1 netRa3 1420.3641638318604
Lbr3 netRa3 netL3 1.2478748845422532e-06
Rbbr3 netL3 node_2 150599.94699341693
Cbr3 netL3 node_2 2.007611429499794e-14

* Branch 4
Rabr4 node_1 netRa4 -6288.153445267598
Lbr4 netRa4 netL4 -1.6984211901391145e-06
Rbbr4 netL4 node_2 -80113.52669092224
Cbr4 netL4 node_2 -1.345066582058904e-14

* Branch 5
Rabr5 node_1 netRa5 -19059.61864984628
Lbr5 netRa5 netL5 -1.0748090317239185e-06
Rbbr5 netL5 node_2 -31974.381807873095
Cbr5 netL5 node_2 -3.2158246530513753e-15

* Branch 6
Rabr6 node_1 netRa6 41171.716014523605
Lbr6 netRa6 netL6 -5.249136740331452e-06
Rbbr6 netL6 node_2 133269.3326801185
Cbr6 netL6 node_2 -8.34764892366965e-16

* Branch 7
Rabr7 node_1 netRa7 -179009.84873316946
Lbr7 netRa7 netL7 2.246106342403787e-05
Rbbr7 netL7 node_2 -597628.5276816767
Cbr7 netL7 node_2 1.974409271007671e-16

* Branch 8
Rabr8 node_1 netRa8 -106.3698467956711
Lbr8 netRa8 netL8 -1.8900705037311493e-07
Rbbr8 netL8 node_2 10713.466699479342
Cbr8 netL8 node_2 -3.342264975024306e-14

* Branch 9
Rabr9 node_1 netRa9 -164688.30836977556
Lbr9 netRa9 netL9 5.4693443889411705e-06
Rbbr9 netL9 node_2 -227439.32835135877
Cbr9 netL9 node_2 1.4203808361899787e-16

* Branch 10
Rabr10 node_1 netRa10 27.11285404881788
Lbr10 netRa10 netL10 -1.3775247808700192e-07
Rbbr10 netL10 node_2 33826.66679001094
Cbr10 netL10 node_2 -2.0405673419146558e-14

* Branch 11
Rabr11 node_1 netRa11 33319.76954778219
Lbr11 netRa11 netL11 1.1900675282283603e-06
Rbbr11 netL11 node_2 66842.20598081908
Cbr11 netL11 node_2 6.853680267811288e-16

* Branch 12
Rabr12 node_1 netRa12 -256817352.30753395
Lbr12 netRa12 netL12 -0.0003666754465629314
Rbbr12 netL12 node_2 -257147791.01212874
Cbr12 netL12 node_2 -5.5602686817779826e-21

* Branch 13
Rabr13 node_1 netRa13 -32.37085881945417
Lbr13 netRa13 netL13 -1.1361908967883745e-07
Rbbr13 netL13 node_2 54862.684585252406
Cbr13 netL13 node_2 -1.3939358263027663e-14

* Branch 14
Rabr14 node_1 netRa14 45884.85290697195
Lbr14 netRa14 netL14 1.4121481676653972e-05
Rbbr14 netL14 node_2 7584689.2477583
Cbr14 netL14 node_2 7.122843326883737e-17

* Branch 15
Rabr15 node_1 netRa15 -25.493103783266765
Lbr15 netRa15 netL15 -1.099482735095784e-07
Rbbr15 netL15 node_2 39039.70924520441
Cbr15 netL15 node_2 -9.204568815385305e-15

* Branch 16
Rabr16 node_1 netRa16 15988.72427187776
Lbr16 netRa16 netL16 1.7084250350420756e-06
Rbbr16 netL16 node_2 323289.9642487844
Cbr16 netL16 node_2 3.91595065279799e-16

* Branch 17
Rabr17 node_1 netRa17 359.0285267867255
Lbr17 netRa17 netL17 -1.3078269828073616e-07
Rbbr17 netL17 node_2 29394.471647759474
Cbr17 netL17 node_2 -5.270388306200524e-15

* Branch 18
Rabr18 node_1 netRa18 -35507.681526097906
Lbr18 netRa18 netL18 -1.7192583396913497e-07
Rbbr18 netL18 node_2 -37207.77962725576
Cbr18 netL18 node_2 -1.7326286293166642e-16

* Branch 19
Rabr19 node_1 netRa19 -171487.47313678602
Lbr19 netRa19 netL19 1.0274714270402394e-05
Rbbr19 netL19 node_2 -1213476.2640570183
Cbr19 netL19 node_2 4.3204311660952656e-17

* Branch 20
Rabr20 node_1 netRa20 10252.049832673332
Lbr20 netRa20 netL20 -1.4438270388838074e-07
Rbbr20 netL20 node_2 14000.768591880498
Cbr20 netL20 node_2 -8.996734958094348e-16

* Branch 21
Rabr21 node_1 netRa21 287.65518298389344
Lbr21 netRa21 netL21 -7.276020156404963e-08
Rbbr21 netL21 node_2 26267.30691942779
Cbr21 netL21 node_2 -5.364492899899159e-15

* Branch 22
Rabr22 node_1 netRa22 -1117.4022519848384
Lbr22 netRa22 netL22 -1.3374866580654672e-07
Rbbr22 netL22 node_2 70649.9470176929
Cbr22 netL22 node_2 -2.9318082773320994e-15

* Branch 23
Rabr23 node_1 netRa23 -176013.7938886835
Lbr23 netRa23 netL23 1.7438700991893275e-06
Rbbr23 netL23 node_2 -228000.4473534987
Cbr23 netL23 node_2 4.0947716439552506e-17

* Branch 24
Rabr24 node_1 netRa24 108.9309860369615
Lbr24 netRa24 netL24 -6.592997137690573e-08
Rbbr24 netL24 node_2 48108.69092786519
Cbr24 netL24 node_2 -4.72824084150829e-15

.ends


* Y'13
.subckt yp13 node_1 node_3
* Branch 0
Rabr0 node_1 netRa0 -1944.9977231079529
Lbr0 netRa0 netL0 -3.2041161848934204e-07
Rbbr0 netL0 node_3 390.1274762941064
Cbr0 netL0 node_3 -4.957170864358547e-13

* Branch 1
Rabr1 node_1 netRa1 -783.5122862386611
Lbr1 netRa1 netL1 1.3913208477095765e-06
Rbbr1 netL1 node_3 -61494.06042191481
Cbr1 netL1 node_3 1.7985264021263132e-14

* Branch 2
Rabr2 node_1 netRa2 4799.378229677052
Lbr2 netRa2 netL2 -5.27601926116265e-06
Rbbr2 netL2 node_3 195210.27029866423
Cbr2 netL2 node_3 -4.683056689860749e-15

* Branch 3
Rabr3 node_1 netRa3 138.38065199000448
Lbr3 netRa3 netL3 -3.542126522543165e-07
Rbbr3 netL3 node_3 11827.625103097425
Cbr3 netL3 node_3 -7.05652614188815e-14

* Branch 4
Rabr4 node_1 netRa4 -1130.4343657608226
Lbr4 netRa4 netL4 -5.324893664143948e-07
Rbbr4 netL4 node_3 31842.552531243167
Cbr4 netL4 node_3 -4.820908158527804e-14

* Branch 5
Rabr5 node_1 netRa5 -38996.66773540508
Lbr5 netRa5 netL5 -1.0946926810186583e-06
Rbbr5 netL5 node_3 -43628.9653777177
Cbr5 netL5 node_3 -8.299820613103469e-16

* Branch 6
Rabr6 node_1 netRa6 -1788.7911453773331
Lbr6 netRa6 netL6 -9.288691852661547e-07
Rbbr6 netL6 node_3 -189502.36070072762
Cbr6 netL6 node_3 -6.76176980510136e-15

* Branch 7
Rabr7 node_1 netRa7 11.885821800483201
Lbr7 netRa7 netL7 -2.1015359187043693e-07
Rbbr7 netL7 node_3 59116.29010817762
Cbr7 netL7 node_3 -3.012007637178824e-14

* Branch 8
Rabr8 node_1 netRa8 3335.953668381816
Lbr8 netRa8 netL8 8.690878320149047e-07
Rbbr8 netL8 node_3 291037.18684668175
Cbr8 netL8 node_3 7.114719401491171e-15

* Branch 9
Rabr9 node_1 netRa9 6579.922552968877
Lbr9 netRa9 netL9 2.6573717014681144e-06
Rbbr9 netL9 node_3 584749.3750098341
Cbr9 netL9 node_3 1.0476541056609114e-15

* Branch 10
Rabr10 node_1 netRa10 -34.59144426051895
Lbr10 netRa10 netL10 -1.3498312262460776e-07
Rbbr10 netL10 node_3 48157.31901102084
Cbr10 netL10 node_3 -2.0855997213799045e-14

* Branch 11
Rabr11 node_1 netRa11 7827.396757057292
Lbr11 netRa11 netL11 1.8347885647849298e-06
Rbbr11 netL11 node_3 -584843.2906716595
Cbr11 netL11 node_3 8.98252750045755e-16

* Branch 12
Rabr12 node_1 netRa12 -6781.897567663409
Lbr12 netRa12 netL12 -1.5290929209266088e-06
Rbbr12 netL12 node_3 -287408.19319189026
Cbr12 netL12 node_3 -1.0131292073993267e-15

* Branch 13
Rabr13 node_1 netRa13 59.9701192826903
Lbr13 netRa13 netL13 -1.2298707765471878e-07
Rbbr13 netL13 node_3 37413.34697516974
Cbr13 netL13 node_3 -1.2849367139784159e-14

* Branch 14
Rabr14 node_1 netRa14 -5035.97778134579
Lbr14 netRa14 netL14 2.0918960198763186e-06
Rbbr14 netL14 node_3 -548212.8062145475
Cbr14 netL14 node_3 4.793149119023644e-16

* Branch 15
Rabr15 node_1 netRa15 142.82641873182018
Lbr15 netRa15 netL15 -1.0298366446489455e-07
Rbbr15 netL15 node_3 23276.756594582544
Cbr15 netL15 node_3 -9.760385552460548e-15

* Branch 16
Rabr16 node_1 netRa16 -63.710395255729445
Lbr16 netRa16 netL16 -9.061361588028837e-08
Rbbr16 netL16 node_3 170081.79708009417
Cbr16 netL16 node_3 -7.770164931037865e-15

* Branch 17
Rabr17 node_1 netRa17 898883.8338594382
Lbr17 netRa17 netL17 8.810470046977881e-06
Rbbr17 netL17 node_3 1027308.9803957336
Cbr17 netL17 node_3 9.901021727723514e-18

* Branch 18
Rabr18 node_1 netRa18 -629512.4230065384
Lbr18 netRa18 netL18 1.1441369497667659e-06
Rbbr18 netL18 node_3 -632429.5155593145
Cbr18 netL18 node_3 2.628248739564418e-18

* Branch 19
Rabr19 node_1 netRa19 -48.1111895958512
Lbr19 netRa19 netL19 -7.552481628613766e-08
Rbbr19 netL19 node_3 83589.16238449015
Cbr19 netL19 node_3 -6.848970548212594e-15

* Branch 20
Rabr20 node_1 netRa20 -2861.652194572852
Lbr20 netRa20 netL20 1.6833005995102363e-07
Rbbr20 netL20 node_3 -16530.686669686304
Cbr20 netL20 node_3 2.3831664802022267e-15

* Branch 21
Rabr21 node_1 netRa21 -34858.310295246825
Lbr21 netRa21 netL21 -3.091790556596975e-06
Rbbr21 netL21 node_3 -998349.6084962044
Cbr21 netL21 node_3 -1.2318557933879589e-16

* Branch 22
Rabr22 node_1 netRa22 1293.1085315362327
Lbr22 netRa22 netL22 -5.3842812997684395e-08
Rbbr22 netL22 node_3 5042.7531397758985
Cbr22 netL22 node_3 -5.330950097235006e-15

* Branch 23
Rabr23 node_1 netRa23 -152656.43798799804
Lbr23 netRa23 netL23 1.4017305323978582e-06
Rbbr23 netL23 node_3 -191548.59612316336
Cbr23 netL23 node_3 4.536346212358475e-17

* Branch 24
Rabr24 node_1 netRa24 161.09072320203816
Lbr24 netRa24 netL24 -6.65116857724143e-08
Rbbr24 netL24 node_3 41368.918117249916
Cbr24 netL24 node_3 -4.679231699136778e-15

.ends


* Y'14
.subckt yp14 node_1 node_4
* Branch 0
Rabr0 node_1 netRa0 -2239.1457042987895
Lbr0 netRa0 netL0 -1.2542625441914261e-06
Rbbr0 netL0 node_4 2759.4378183652825
Cbr0 netL0 node_4 -3.832449138885801e-14

* Branch 1
Rabr1 node_1 netRa1 53127.656909406636
Lbr1 netRa1 netL1 -7.960534896222015e-06
Rbbr1 netL1 node_4 97899.72804992906
Cbr1 netL1 node_4 -1.456118017788345e-15

* Branch 2
Rabr2 node_1 netRa2 -196667.66480880827
Lbr2 netRa2 netL2 2.7123418756508443e-05
Rbbr2 netL2 node_4 -340684.50650977955
Cbr2 netL2 node_4 3.947872630842864e-16

* Branch 3
Rabr3 node_1 netRa3 -19498.23749175193
Lbr3 netRa3 netL3 3.5588080565180353e-06
Rbbr3 netL3 node_4 -41882.359884363104
Cbr3 netL3 node_4 3.7981358696879935e-15

* Branch 4
Rabr4 node_1 netRa4 1514.2135336943402
Lbr4 netRa4 netL4 -4.737389098657475e-07
Rbbr4 netL4 node_4 4714.788376470156
Cbr4 netL4 node_4 -3.552352940671879e-14

* Branch 5
Rabr5 node_1 netRa5 38275.51666050238
Lbr5 netRa5 netL5 9.981504483989647e-07
Rbbr5 netL5 node_4 42120.183303969396
Cbr5 netL5 node_4 7.825494831203662e-16

* Branch 6
Rabr6 node_1 netRa6 94.72970548410542
Lbr6 netRa6 netL6 2.399950249661017e-06
Rbbr6 netL6 node_4 -342166.2496461066
Cbr6 netL6 node_4 2.6427243944340586e-15

* Branch 7
Rabr7 node_1 netRa7 14671.339288725088
Lbr7 netRa7 netL7 -1.1157441575292214e-05
Rbbr7 netL7 node_4 982982.3256951151
Cbr7 netL7 node_4 -5.589651634195936e-16

* Branch 8
Rabr8 node_1 netRa8 8.78021296119484
Lbr8 netRa8 netL8 -1.767435955445205e-07
Rbbr8 netL8 node_4 8306.790979990998
Cbr8 netL8 node_4 -3.535291524812065e-14

* Branch 9
Rabr9 node_1 netRa9 60775.78694920969
Lbr9 netRa9 netL9 -6.4693953188323424e-06
Rbbr9 netL9 node_4 285194.5148165868
Cbr9 netL9 node_4 -3.424830537871665e-16

* Branch 10
Rabr10 node_1 netRa10 -28880.852413511184
Lbr10 netRa10 netL10 3.5085028653026682e-06
Rbbr10 netL10 node_4 -160388.34959628826
Cbr10 netL10 node_4 6.574374616051664e-16

* Branch 11
Rabr11 node_1 netRa11 -8928984.079137525
Lbr11 netRa11 netL11 1.4626555320084862e-05
Rbbr11 netL11 node_4 -8943569.006327514
Cbr11 netL11 node_4 1.8132679658128031e-19

* Branch 12
Rabr12 node_1 netRa12 -798472.6839694602
Lbr12 netRa12 netL12 -1.2664252602158528e-05
Rbbr12 netL12 node_4 -927113.7610243417
Cbr12 netL12 node_4 -1.7383473920434963e-17

* Branch 13
Rabr13 node_1 netRa13 124955.92168986655
Lbr13 netRa13 netL13 3.376205073285995e-06
Rbbr13 netL13 node_4 185179.1371902112
Cbr13 netL13 node_4 1.524687986396753e-16

* Branch 14
Rabr14 node_1 netRa14 -10471.774250429182
Lbr14 netRa14 netL14 3.5309514441981555e-06
Rbbr14 netL14 node_4 -810009.0236068285
Cbr14 netL14 node_4 2.8289552323598453e-16

* Branch 15
Rabr15 node_1 netRa15 3803.1580656215738
Lbr15 netRa15 netL15 -1.1818339080016357e-06
Rbbr15 netL15 node_4 191289.5692419299
Cbr15 netL15 node_4 -8.387459189170141e-16

* Branch 16
Rabr16 node_1 netRa16 -1246038.2191419695
Lbr16 netRa16 netL16 1.778976021831119e-05
Rbbr16 netL16 node_4 -1599538.3056978947
Cbr16 netL16 node_4 8.743510437949534e-18

* Branch 17
Rabr17 node_1 netRa17 135947.41552386712
Lbr17 netRa17 netL17 2.7341108631828654e-06
Rbbr17 netL17 node_4 221101.47409435574
Cbr17 netL17 node_4 9.829415662028323e-17

* Branch 18
Rabr18 node_1 netRa18 -208.367109446998
Lbr18 netRa18 netL18 -9.892804436877077e-09
Rbbr18 netL18 node_4 291.62991089009
Cbr18 netL18 node_4 -1.1298539937028145e-13

* Branch 19
Rabr19 node_1 netRa19 -1829875.5420123434
Lbr19 netRa19 netL19 -1.910264606072896e-05
Rbbr19 netL19 node_4 -2225464.775006587
Cbr19 netL19 node_4 -4.810556185283772e-18

* Branch 20
Rabr20 node_1 netRa20 406.64074531739436
Lbr20 netRa20 netL20 3.6106518675566133e-07
Rbbr20 netL20 node_4 -102145.8743762264
Cbr20 netL20 node_4 1.3489907888306016e-15

* Branch 21
Rabr21 node_1 netRa21 389.7674255080684
Lbr21 netRa21 netL21 1.390131381158539e-06
Rbbr21 netL21 node_4 -1230032.532153505
Cbr21 netL21 node_4 2.839792057795709e-16

* Branch 22
Rabr22 node_1 netRa22 180721.47029478033
Lbr22 netRa22 netL22 -8.545816432297297e-07
Rbbr22 netL22 node_4 190575.76810292088
Cbr22 netL22 node_4 -2.3356857126737213e-17

* Branch 23
Rabr23 node_1 netRa23 -86882.06570860188
Lbr23 netRa23 netL23 1.1167906054756378e-06
Rbbr23 netL23 node_4 -129347.62012454636
Cbr23 netL23 node_4 9.206493692744433e-17

* Branch 24
Rabr24 node_1 netRa24 -3104.597315228933
Lbr24 netRa24 netL24 7.541127934084467e-07
Rbbr24 netL24 node_4 -354900.5765629499
Cbr24 netL24 node_4 4.1069064420184607e-16

.ends


* Y'22
.subckt yp22 node_2 node_ref
* Branch 0
Rabr0 node_2 netRa0 11899.825265252772
Lbr0 netRa0 netL0 -9.356753175084473e-07
Rbbr0 netL0 node_ref 13371.51886552739
Cbr0 netL0 node_ref -3.1214041157076246e-15

* Branch 1
Rabr1 node_2 netRa1 39.410438209014245
Lbr1 netRa1 netL1 1.6829328214043804e-07
Rbbr1 netL1 node_ref -62101.76240435409
Cbr1 netL1 node_ref 1.507029892054777e-13

* Branch 2
Rabr2 node_2 netRa2 1447.465878698852
Lbr2 netRa2 netL2 2.1286086783522134e-06
Rbbr2 netL2 node_ref 170940.65683528795
Cbr2 netL2 node_ref 1.1799340166528538e-14

* Branch 3
Rabr3 node_2 netRa3 52.96358985937849
Lbr3 netRa3 netL3 2.3756893828328224e-07
Rbbr3 netL3 node_ref -16016.796911076586
Cbr3 netL3 node_ref 1.0680958130973997e-13

* Branch 4
Rabr4 node_2 netRa4 444.02672863761546
Lbr4 netRa4 netL4 -9.307934027228115e-07
Rbbr4 netL4 node_ref 11991.715934747876
Cbr4 netL4 node_ref -2.5647783533200213e-14

* Branch 5
Rabr5 node_2 netRa5 -961.6778464599976
Lbr5 netRa5 netL5 -2.839810058012946e-07
Rbbr5 netL5 node_ref 6219.403466592227
Cbr5 netL5 node_ref -3.479294558753787e-14

* Branch 6
Rabr6 node_2 netRa6 131.67641569906064
Lbr6 netRa6 netL6 1.3527198042711046e-07
Rbbr6 netL6 node_ref -123947.46349023197
Cbr6 netL6 node_ref 4.6923151832585305e-14

* Branch 7
Rabr7 node_2 netRa7 648.6499415440188
Lbr7 netRa7 netL7 6.248483896422913e-07
Rbbr7 netL7 node_ref 185804.3439410934
Cbr7 netL7 node_ref 1.0096870063408314e-14

* Branch 8
Rabr8 node_2 netRa8 -54.312065335111036
Lbr8 netRa8 netL8 1.273217480437132e-07
Rbbr8 netL8 node_ref -5436.302254769953
Cbr8 netL8 node_ref 4.863679184043468e-14

* Branch 9
Rabr9 node_2 netRa9 256.8755078000526
Lbr9 netRa9 netL9 1.0111010946674652e-07
Rbbr9 netL9 node_ref 21420.004785970323
Cbr9 netL9 node_ref 2.7513800898914305e-14

* Branch 10
Rabr10 node_2 netRa10 -96.78774742946035
Lbr10 netRa10 netL10 8.69053636178253e-08
Rbbr10 netL10 node_ref -13155.528186824262
Cbr10 netL10 node_ref 3.2132536383149157e-14

* Branch 11
Rabr11 node_2 netRa11 568.2519704353991
Lbr11 netRa11 netL11 6.869624343323127e-08
Rbbr11 netL11 node_ref 20660.37709175002
Cbr11 netL11 node_ref 2.3023178744148987e-14

* Branch 12
Rabr12 node_2 netRa12 -346012.5996379677
Lbr12 netRa12 netL12 1.2647856928448895e-05
Rbbr12 netL12 node_ref -627116.0644147012
Cbr12 netL12 node_ref 5.623035468198689e-17

* Branch 13
Rabr13 node_2 netRa13 171.66755662529042
Lbr13 netRa13 netL13 1.1391824172612303e-07
Rbbr13 netL13 node_ref -840742.5868701027
Cbr13 netL13 node_ref 1.3897391978642377e-14

* Branch 14
Rabr14 node_2 netRa14 -3727.4410407487835
Lbr14 netRa14 netL14 8.673251250411329e-07
Rbbr14 netL14 node_ref -154197.3410183908
Cbr14 netL14 node_ref 1.1385701551398566e-15

* Branch 15
Rabr15 node_2 netRa15 51.57100437326929
Lbr15 netRa15 netL15 4.768316948630017e-08
Rbbr15 netL15 node_ref -24336.882068985087
Cbr15 netL15 node_ref 2.1255071055575427e-14

* Branch 16
Rabr16 node_2 netRa16 -162.62876919458031
Lbr16 netRa16 netL16 2.2277989771827553e-07
Rbbr16 netL16 node_ref -144711.65136837514
Cbr16 netL16 node_ref 3.1557072496873297e-15

* Branch 17
Rabr17 node_2 netRa17 -235.81936066272684
Lbr17 netRa17 netL17 5.1634021722118955e-08
Rbbr17 netL17 node_ref -9175.902664504918
Cbr17 netL17 node_ref 1.3167002611120543e-14

* Branch 18
Rabr18 node_2 netRa18 784.6159694518238
Lbr18 netRa18 netL18 2.3648446504896518e-08
Rbbr18 netL18 node_ref -1204.8302784032971
Cbr18 netL18 node_ref 4.5520824288647154e-14

* Branch 19
Rabr19 node_2 netRa19 -39660.66888869082
Lbr19 netRa19 netL19 1.6169208527172916e-06
Rbbr19 netL19 node_ref -155878.6703941045
Cbr19 netL19 node_ref 2.3837627595648534e-16

* Branch 20
Rabr20 node_2 netRa20 -2112.4177486860226
Lbr20 netRa20 netL20 3.5242651412254414e-08
Rbbr20 netL20 node_ref -3175.6656682224298
Cbr20 netL20 node_ref 4.608932084347539e-15

* Branch 21
Rabr21 node_2 netRa21 -140.43023077590942
Lbr21 netRa21 netL21 3.451017127801105e-08
Rbbr21 netL21 node_ref -12264.789022399043
Cbr21 netL21 node_ref 1.1304630589227952e-14

* Branch 22
Rabr22 node_2 netRa22 267.00814142301533
Lbr22 netRa22 netL22 1.1204022129089394e-08
Rbbr22 netL22 node_ref 2992.5326184258947
Cbr22 netL22 node_ref 3.137958499286269e-14

* Branch 23
Rabr23 node_2 netRa23 3744.917844311574
Lbr23 netRa23 netL23 7.913075236135758e-08
Rbbr23 netL23 node_ref 9885.577492080047
Cbr23 netL23 node_ref 2.4584158261524104e-15

* Branch 24
Rabr24 node_2 netRa24 -386.9334966930026
Lbr24 netRa24 netL24 7.203164757615866e-08
Rbbr24 netL24 node_ref -28794.309211489526
Cbr24 netL24 node_ref 4.2792538902186915e-15

.ends


* Y'23
.subckt yp23 node_2 node_3
* Branch 0
Rabr0 node_2 netRa0 1878.7434463350305
Lbr0 netRa0 netL0 2.716050062809983e-07
Rbbr0 netL0 node_3 -488.3721211833202
Cbr0 netL0 node_3 4.735538139222589e-13

* Branch 1
Rabr1 node_2 netRa1 -566.1231343658915
Lbr1 netRa1 netL1 -2.716804833250842e-06
Rbbr1 netL1 node_3 807491.0570484446
Cbr1 netL1 node_3 -9.335961622173844e-15

* Branch 2
Rabr2 node_2 netRa2 -2069.9372527546066
Lbr2 netRa2 netL2 1.3193243558644743e-05
Rbbr2 netL2 node_3 -1528967.9830714974
Cbr2 netL2 node_3 1.917373543597776e-15

* Branch 3
Rabr3 node_2 netRa3 -218.54454799741364
Lbr3 netRa3 netL3 -2.950123599858149e-07
Rbbr3 netL3 node_3 174712.49724486456
Cbr3 netL3 node_3 -8.583587399421669e-14

* Branch 4
Rabr4 node_2 netRa4 4139.08671273094
Lbr4 netRa4 netL4 1.3899473954742522e-06
Rbbr4 netL4 node_3 279618.7006991199
Cbr4 netL4 node_3 1.757171981662707e-14

* Branch 5
Rabr5 node_2 netRa5 11274.147604235575
Lbr5 netRa5 netL5 4.5654304835822027e-07
Rbbr5 netL5 node_3 14471.319590007204
Cbr5 netL5 node_3 4.141097995469134e-15

* Branch 6
Rabr6 node_2 netRa6 -525.4267652117371
Lbr6 netRa6 netL6 -4.089103481692751e-07
Rbbr6 netL6 node_3 -462541.00523723563
Cbr6 netL6 node_3 -1.5488600282180154e-14

* Branch 7
Rabr7 node_2 netRa7 -1469.0122301039455
Lbr7 netRa7 netL7 3.1868946971049534e-06
Rbbr7 netL7 node_3 -522551.41504366515
Cbr7 netL7 node_3 1.9810246460219227e-15

* Branch 8
Rabr8 node_2 netRa8 -299.3087830585994
Lbr8 netRa8 netL8 -1.8670181245886195e-07
Rbbr8 netL8 node_3 16733.771832914696
Cbr8 netL8 node_3 -3.410193571116368e-14

* Branch 9
Rabr9 node_2 netRa9 -370.32509095554275
Lbr9 netRa9 netL9 -1.366905632430185e-07
Rbbr9 netL9 node_3 -26393.853060035774
Cbr9 netL9 node_3 -2.0309989302502512e-14

* Branch 10
Rabr10 node_2 netRa10 274977.3206391912
Lbr10 netRa10 netL10 3.941854906433503e-06
Rbbr10 netL10 node_3 295430.9619592617
Cbr10 netL10 node_3 4.9409741450645546e-17

* Branch 11
Rabr11 node_2 netRa11 -2486.205321053006
Lbr11 netRa11 netL11 -1.5684365087315896e-07
Rbbr11 netL11 node_3 -12447.095046843466
Cbr11 netL11 node_3 -8.298007585061867e-15

* Branch 12
Rabr12 node_2 netRa12 -5452.6913894195595
Lbr12 netRa12 netL12 2.0020175950404344e-06
Rbbr12 netL12 node_3 -344237.2962683014
Cbr12 netL12 node_3 7.799510539360693e-16

* Branch 13
Rabr13 node_2 netRa13 2415.6287531707003
Lbr13 netRa13 netL13 -8.194435485853172e-07
Rbbr13 netL13 node_3 116436.90038449822
Cbr13 netL13 node_3 -1.8915338457242704e-15

* Branch 14
Rabr14 node_2 netRa14 81813.31143319391
Lbr14 netRa14 netL14 4.1390597160132915e-06
Rbbr14 netL14 node_3 304489.51800844114
Cbr14 netL14 node_3 1.7880050903045977e-16

* Branch 15
Rabr15 node_2 netRa15 -11012.156875207103
Lbr15 netRa15 netL15 -8.226728389547287e-07
Rbbr15 netL15 node_3 -89444.19016703242
Cbr15 netL15 node_3 -1.0780093756037102e-15

* Branch 16
Rabr16 node_2 netRa16 -48220.181331973385
Lbr16 netRa16 netL16 3.3221669771452705e-06
Rbbr16 netL16 node_3 -343704.42363435996
Cbr16 netL16 node_3 1.8213306441038093e-16

* Branch 17
Rabr17 node_2 netRa17 6118.119679345853
Lbr17 netRa17 netL17 -4.1165967509997705e-07
Rbbr17 netL17 node_3 37883.53771026322
Cbr17 netL17 node_3 -1.4213329593132465e-15

* Branch 18
Rabr18 node_2 netRa18 -3025.0160593983114
Lbr18 netRa18 netL18 -4.1672986399766405e-08
Rbbr18 netL18 node_3 -6043.350887408087
Cbr18 netL18 node_3 -7.813423739879718e-15

* Branch 19
Rabr19 node_2 netRa19 -890084.3429760338
Lbr19 netRa19 netL19 -7.178409940060014e-06
Rbbr19 netL19 node_3 -1004264.521040274
Cbr19 netL19 node_3 -8.18802994266091e-18

* Branch 20
Rabr20 node_2 netRa20 11669.405224452785
Lbr20 netRa20 netL20 1.5572621869285582e-07
Rbbr20 netL20 node_3 16492.567222791473
Cbr20 netL20 node_3 9.110683568887242e-16

* Branch 21
Rabr21 node_2 netRa21 -113.22927861799278
Lbr21 netRa21 netL21 -4.292548459127856e-07
Rbbr21 netL21 node_3 377635.0446639533
Cbr21 netL21 node_3 -9.196440888949792e-16

* Branch 22
Rabr22 node_2 netRa22 214.54090819101035
Lbr22 netRa22 netL22 -2.352671839883079e-08
Rbbr22 netL22 node_3 2947.417406215836
Cbr22 netL22 node_3 -1.5213423934007224e-14

* Branch 23
Rabr23 node_2 netRa23 -3813.341596602461
Lbr23 netRa23 netL23 -1.197308881415041e-07
Rbbr23 netL23 node_3 -18706.122837048504
Cbr23 netL23 node_3 -2.0824447138604757e-15

* Branch 24
Rabr24 node_2 netRa24 210242.27845173224
Lbr24 netRa24 netL24 3.0533218823970747e-06
Rbbr24 netL24 node_3 358057.5301587007
Cbr24 netL24 node_3 4.224358785845284e-17

.ends


* Y'24
.subckt yp24 node_2 node_4
* Branch 0
Rabr0 node_2 netRa0 -2546.267756488449
Lbr0 netRa0 netL0 -2.2912484106604106e-07
Rbbr0 netL0 node_4 64848.82576637552
Cbr0 netL0 node_4 -1.2036286007754727e-13

* Branch 1
Rabr1 node_2 netRa1 -318662.26685069833
Lbr1 netRa1 netL1 2.5842154203584815e-05
Rbbr1 netL1 node_4 -399119.66118222947
Cbr1 netL1 node_4 1.977184759414624e-16

* Branch 2
Rabr2 node_2 netRa2 1275204.6387086713
Lbr2 netRa2 netL2 -9.154214813166323e-05
Rbbr2 netL2 node_4 1531245.9784114202
Cbr2 netL2 node_4 -4.626906175780469e-17

* Branch 3
Rabr3 node_2 netRa3 292594.13263425423
Lbr3 netRa3 netL3 -1.862870878903398e-05
Rbbr3 netL3 node_4 337196.8789510712
Cbr3 netL3 node_4 -1.7958143370246584e-16

* Branch 4
Rabr4 node_2 netRa4 -52648.353751984185
Lbr4 netRa4 netL4 4.771890989131235e-06
Rbbr4 netL4 node_4 -66589.23922603535
Cbr4 netL4 node_4 1.0876400064546627e-15

* Branch 5
Rabr5 node_2 netRa5 -738549.962122701
Lbr5 netRa5 netL5 5.664193708637837e-06
Rbbr5 netL5 node_4 -743332.6527647702
Cbr5 netL5 node_4 9.720539297102382e-18

* Branch 6
Rabr6 node_2 netRa6 -46487.303681485144
Lbr6 netRa6 netL6 -1.1504788611737104e-05
Rbbr6 netL6 node_4 -673167.9518509267
Cbr6 netL6 node_4 -5.130717492637134e-16

* Branch 7
Rabr7 node_2 netRa7 160652.17530993558
Lbr7 netRa7 netL7 4.793586986623393e-05
Rbbr7 netL7 node_4 2820722.5763619384
Cbr7 netL7 node_4 1.245524735315404e-16

* Branch 8
Rabr8 node_2 netRa8 6506.685185255346
Lbr8 netRa8 netL8 2.52016646579372e-06
Rbbr8 netL8 node_4 -514265.1767546822
Cbr8 netL8 node_4 2.5133870405289132e-15

* Branch 9
Rabr9 node_2 netRa9 -105793.83534434467
Lbr9 netRa9 netL9 3.138702498053051e-05
Rbbr9 netL9 node_4 -2750830.889036701
Cbr9 netL9 node_4 8.625863161838073e-17

* Branch 10
Rabr10 node_2 netRa10 245949.0564895827
Lbr10 netRa10 netL10 -3.325205988476962e-05
Rbbr10 netL10 node_4 1612680.3740404944
Cbr10 netL10 node_4 -7.169929411588324e-17

* Branch 11
Rabr11 node_2 netRa11 593810.5437448255
Lbr11 netRa11 netL11 8.701707030525105e-06
Rbbr11 netL11 node_4 680010.033959373
Cbr11 netL11 node_4 2.369166390760842e-17

* Branch 12
Rabr12 node_2 netRa12 200795.20680653647
Lbr12 netRa12 netL12 1.5560215324470904e-05
Rbbr12 netL12 node_4 1024693.6757937033
Cbr12 netL12 node_4 8.198483594705421e-17

* Branch 13
Rabr13 node_2 netRa13 -405524.1148036446
Lbr13 netRa13 netL13 -1.632275374736032e-05
Rbbr13 netL13 node_4 -849033.8016558954
Cbr13 netL13 node_4 -5.065503422096245e-17

* Branch 14
Rabr14 node_2 netRa14 552757.7958283821
Lbr14 netRa14 netL14 4.272261457666584e-05
Rbbr14 netL14 node_4 4211085.713015685
Cbr14 netL14 node_4 2.0577836034282714e-17

* Branch 15
Rabr15 node_2 netRa15 -36257.99134800006
Lbr15 netRa15 netL15 7.93730624776622e-06
Rbbr15 netL15 node_4 -1071250.7002411722
Cbr15 netL15 node_4 1.2310661610836169e-16

* Branch 16
Rabr16 node_2 netRa16 97627.50169601613
Lbr16 netRa16 netL16 7.326951713331706e-06
Rbbr16 netL16 node_4 975046.5970862678
Cbr16 netL16 node_4 8.644092969866185e-17

* Branch 17
Rabr17 node_2 netRa17 -217256.85502824173
Lbr17 netRa17 netL17 -5.2660491706874624e-06
Rbbr17 netL17 node_4 -418252.24216924835
Cbr17 netL17 node_4 -6.367852716980416e-17

* Branch 18
Rabr18 node_2 netRa18 -573.4571864610789
Lbr18 netRa18 netL18 -1.3693467204993366e-08
Rbbr18 netL18 node_4 1629.7653008663467
Cbr18 netL18 node_4 -6.43615153037002e-14

* Branch 19
Rabr19 node_2 netRa19 44999.53374825674
Lbr19 netRa19 netL19 7.258552440918095e-06
Rbbr19 netL19 node_4 3724619.2682685233
Cbr19 netL19 node_4 7.036166654211707e-17

* Branch 20
Rabr20 node_2 netRa20 22717.139514520666
Lbr20 netRa20 netL20 -5.53383969828434e-07
Rbbr20 netL20 node_4 45791.25406100634
Cbr20 netL20 node_4 -4.417586350493583e-16

* Branch 21
Rabr21 node_2 netRa21 19619.40760396194
Lbr21 netRa21 netL21 9.503291245782621e-07
Rbbr21 netL21 node_4 157210.59422473906
Cbr21 netL21 node_4 3.6344572062897606e-16

* Branch 22
Rabr22 node_2 netRa22 -4387.772003139615
Lbr22 netRa22 netL22 -9.375874809536421e-08
Rbbr22 netL22 node_4 -11613.026665083296
Cbr22 netL22 node_4 -2.5615680372351e-15

* Branch 23
Rabr23 node_2 netRa23 -5313143.151615969
Lbr23 netRa23 netL23 -5.163557359935968e-06
Rbbr23 netL23 node_4 -5329263.497156545
Cbr23 netL23 node_4 -1.8346186460125907e-19

* Branch 24
Rabr24 node_2 netRa24 6583.39144832567
Lbr24 netRa24 netL24 7.203262704276304e-07
Rbbr24 netL24 node_4 367069.67927760916
Cbr24 netL24 node_4 4.2596894167965816e-16

.ends


* Y'33
.subckt yp33 node_3 node_ref
* Branch 0
Rabr0 node_3 netRa0 -958.8191953802551
Lbr0 netRa0 netL0 -1.6775820317396718e-07
Rbbr0 netL0 node_ref 185.2756326000121
Cbr0 netL0 node_ref -9.767838348014351e-13

* Branch 1
Rabr1 node_3 netRa1 10602.507269717235
Lbr1 netRa1 netL1 -6.256699732877323e-06
Rbbr1 netL1 node_ref 131868.0037863145
Cbr1 netL1 node_ref -3.725337557298574e-15

* Branch 2
Rabr2 node_3 netRa2 -25839.52356675218
Lbr2 netRa2 netL2 1.77251411925703e-05
Rbbr2 netL2 node_ref -451995.2136593348
Cbr2 netL2 node_ref 1.3473840900302953e-15

* Branch 3
Rabr3 node_3 netRa3 52.47339046047397
Lbr3 netRa3 netL3 1.7152648738426242e-07
Rbbr3 netL3 node_ref -13469.573773130835
Cbr3 netL3 node_ref 1.480210679410423e-13

* Branch 4
Rabr4 node_3 netRa4 308.3342687833435
Lbr4 netRa4 netL4 1.6032478637373285e-07
Rbbr4 netL4 node_ref -7289.663335869944
Cbr4 netL4 node_ref 1.611685847819906e-13

* Branch 5
Rabr5 node_3 netRa5 -1433.9582865529158
Lbr5 netRa5 netL5 -1.6111709902628384e-07
Rbbr5 netL5 node_ref -22531.3785415364
Cbr5 netL5 node_ref -4.9732390401055545e-14

* Branch 6
Rabr6 node_3 netRa6 484.43853426133705
Lbr6 netRa6 netL6 2.6902426039597637e-07
Rbbr6 netL6 node_ref 65224.65001277617
Cbr6 netL6 node_ref 2.3394017140885207e-14

* Branch 7
Rabr7 node_3 netRa7 -18.073547620493482
Lbr7 netRa7 netL7 2.2747186226748032e-07
Rbbr7 netL7 node_ref -61487.12208141491
Cbr7 netL7 node_ref 2.78243389176025e-14

* Branch 8
Rabr8 node_3 netRa8 -495.09661722873375
Lbr8 netRa8 netL8 2.8534457180424746e-07
Rbbr8 netL8 node_ref -9456.43164593266
Cbr8 netL8 node_ref 2.0773229430095553e-14

* Branch 9
Rabr9 node_3 netRa9 533.613101487063
Lbr9 netRa9 netL9 1.5323548210003315e-07
Rbbr9 netL9 node_ref 21159.316520163164
Cbr9 netL9 node_ref 1.7911528311796836e-14

* Branch 10
Rabr10 node_3 netRa10 -358.53005420482987
Lbr10 netRa10 netL10 1.2710393895017378e-07
Rbbr10 netL10 node_ref -11452.331002997335
Cbr10 netL10 node_ref 2.144006297112123e-14

* Branch 11
Rabr11 node_3 netRa11 3897.6401381437217
Lbr11 netRa11 netL11 3.7337189500355183e-07
Rbbr11 netL11 node_ref 57670.7909673893
Cbr11 netL11 node_ref 4.061426487129371e-15

* Branch 12
Rabr12 node_3 netRa12 -6359.676676852775
Lbr12 netRa12 netL12 -3.45225982301048e-06
Rbbr12 netL12 node_ref -2592936.358346268
Cbr12 netL12 node_ref -4.584579636443494e-16

* Branch 13
Rabr13 node_3 netRa13 12.962136462711603
Lbr13 netRa13 netL13 9.652506818940932e-08
Rbbr13 netL13 node_ref -41806.14092691162
Cbr13 netL13 node_ref 1.6403345375258765e-14

* Branch 14
Rabr14 node_3 netRa14 -34284.662888530125
Lbr14 netRa14 netL14 -2.144131170923503e-06
Rbbr14 netL14 node_ref -179487.7799754724
Cbr14 netL14 node_ref -3.8182000462196297e-16

* Branch 15
Rabr15 node_3 netRa15 156.68106016224633
Lbr15 netRa15 netL15 9.975719411320912e-08
Rbbr15 netL15 node_ref -68146.53533059469
Cbr15 netL15 node_ref 1.0161586272897612e-14

* Branch 16
Rabr16 node_3 netRa16 43.69148314811576
Lbr16 netRa16 netL16 9.401474248009666e-08
Rbbr16 netL16 node_ref -134198.95248834026
Cbr16 netL16 node_ref 7.48870043771915e-15

* Branch 17
Rabr17 node_3 netRa17 -1712.411294972801
Lbr17 netRa17 netL17 3.372926334388979e-07
Rbbr17 netL17 node_ref -56724.0037658875
Cbr17 netL17 node_ref 2.0063679926554126e-15

* Branch 18
Rabr18 node_3 netRa18 73.18733148099174
Lbr18 netRa18 netL18 5.21025859753257e-09
Rbbr18 netL18 node_ref -140.7025293842182
Cbr18 netL18 node_ref 1.9021090514862885e-13

* Branch 19
Rabr19 node_3 netRa19 97.68137551946933
Lbr19 netRa19 netL19 7.582211136344285e-08
Rbbr19 netL19 node_ref -133788.77584173085
Cbr19 netL19 node_ref 6.823169788849299e-15

* Branch 20
Rabr20 node_3 netRa20 -8673.075282303169
Lbr20 netRa20 netL20 -1.4533667653222936e-07
Rbbr20 netL20 node_ref -14513.627016156908
Cbr20 netL20 node_ref -1.3432962659216008e-15

* Branch 21
Rabr21 node_3 netRa21 -2652.485818485537
Lbr21 netRa21 netL21 3.8635879728821493e-07
Rbbr21 netL21 node_ref -100469.46706122464
Cbr21 netL21 node_ref 9.944756270882108e-16

* Branch 22
Rabr22 node_3 netRa22 -21.53396411483869
Lbr22 netRa22 netL22 1.4443142960335439e-08
Rbbr22 netL22 node_ref -2571.442706011755
Cbr22 netL22 node_ref 2.6503060949593746e-14

* Branch 23
Rabr23 node_3 netRa23 11384.781080203633
Lbr23 netRa23 netL23 1.6052493935892715e-07
Rbbr23 netL23 node_ref 19301.693932596645
Cbr23 netL23 node_ref 8.002129605497509e-16

* Branch 24
Rabr24 node_3 netRa24 -333.0175032765135
Lbr24 netRa24 netL24 6.734916071313479e-08
Rbbr24 netL24 node_ref -28369.090739033323
Cbr24 netL24 node_ref 4.584653655644895e-15

.ends


* Y'34
.subckt yp34 node_3 node_4
* Branch 0
Rabr0 node_3 netRa0 1580.9834323363305
Lbr0 netRa0 netL0 4.3437878185109646e-07
Rbbr0 netL0 node_4 -572.449837252497
Cbr0 netL0 node_4 2.2980733748299033e-13

* Branch 1
Rabr1 node_3 netRa1 1725.0054203831512
Lbr1 netRa1 netL1 -5.4739830582107865e-06
Rbbr1 netL1 node_4 330867.4069442054
Cbr1 netL1 node_4 -4.606165342577682e-15

* Branch 2
Rabr2 node_3 netRa2 -11295.578125615366
Lbr2 netRa2 netL2 1.8051380141785326e-05
Rbbr2 netL2 node_4 -891125.660506652
Cbr2 netL2 node_4 1.385466750710835e-15

* Branch 3
Rabr3 node_3 netRa3 -56.46332891573146
Lbr3 netRa3 netL3 2.8260529728849195e-06
Rbbr3 netL3 node_4 -135098.0484177621
Cbr3 netL3 node_4 8.945493149355606e-15

* Branch 4
Rabr4 node_3 netRa4 -974.2275396399424
Lbr4 netRa4 netL4 -4.644749566486492e-07
Rbbr4 netL4 node_4 26706.044565870627
Cbr4 netL4 node_4 -5.532072514547899e-14

* Branch 5
Rabr5 node_3 netRa5 15913.153835219038
Lbr5 netRa5 netL5 1.0005561569248435e-06
Rbbr5 netL5 node_4 30719.911604097713
Cbr5 netL5 node_4 4.122284098805583e-15

* Branch 6
Rabr6 node_3 netRa6 93590.10090209305
Lbr6 netRa6 netL6 -1.1389434366843897e-05
Rbbr6 netL6 node_4 285443.8403497859
Cbr6 netL6 node_4 -3.7418065433061477e-16

* Branch 7
Rabr7 node_3 netRa7 -561077.7133540761
Lbr7 netRa7 netL7 4.828087583579853e-05
Rbbr7 netL7 node_4 -1189962.672921523
Cbr7 netL7 node_4 6.930154920151067e-17

* Branch 8
Rabr8 node_3 netRa8 -778.1795918429192
Lbr8 netRa8 netL8 3.417267012359425e-06
Rbbr8 netL8 node_4 -153245.10016079995
Cbr8 netL8 node_4 1.8211189924561434e-15

* Branch 9
Rabr9 node_3 netRa9 -151382.22119269954
Lbr9 netRa9 netL9 6.053491285111825e-06
Rbbr9 netL9 node_4 -234547.2452358468
Cbr9 netL9 node_4 1.6492606941290962e-16

* Branch 10
Rabr10 node_3 netRa10 87685.33898196211
Lbr10 netRa10 netL10 -3.5457408255918816e-06
Rbbr10 netL10 node_4 136196.4433069433
Cbr10 netL10 node_4 -2.8259664112571527e-16

* Branch 11
Rabr11 node_3 netRa11 2184.282182236759
Lbr11 netRa11 netL11 4.0646181212305696e-07
Rbbr11 netL11 node_4 -311890.1393344307
Cbr11 netL11 node_4 4.029227775965818e-15

* Branch 12
Rabr12 node_3 netRa12 -8633.126245827536
Lbr12 netRa12 netL12 3.6655770866389536e-06
Rbbr12 netL12 node_4 -697018.5751688533
Cbr12 netL12 node_4 4.2747868729595204e-16

* Branch 13
Rabr13 node_3 netRa13 7054.990050875368
Lbr13 netRa13 netL13 -1.6740565215665868e-06
Rbbr13 netL13 node_4 189189.8306492849
Cbr13 netL13 node_4 -9.102549243218514e-16

* Branch 14
Rabr14 node_3 netRa14 503148.8200203598
Lbr14 netRa14 netL14 -1.196774442594707e-05
Rbbr14 netL14 node_4 775387.5515525737
Cbr14 netL14 node_4 -2.968846595693916e-17

* Branch 15
Rabr15 node_3 netRa15 -158109.70517945883
Lbr15 netRa15 netL15 3.574966928009588e-06
Rbbr15 netL15 node_4 -232933.36142236876
Cbr15 netL15 node_4 9.087481987450208e-17

* Branch 16
Rabr16 node_3 netRa16 471678.1955198989
Lbr16 netRa16 netL16 1.4560894263583638e-05
Rbbr16 netL16 node_4 1140476.1934338803
Cbr16 netL16 node_4 2.8345344512983113e-17

* Branch 17
Rabr17 node_3 netRa17 -58792.57335213814
Lbr17 netRa17 netL17 -2.6268963970042103e-06
Rbbr17 netL17 node_4 -260414.75612479454
Cbr17 netL17 node_4 -2.0566476096252923e-16

* Branch 18
Rabr18 node_3 netRa18 -24.527294165670455
Lbr18 netRa18 netL18 -1.1807405122060127e-08
Rbbr18 netL18 node_4 342.5851682590788
Cbr18 netL18 node_4 -5.916740257580977e-14

* Branch 19
Rabr19 node_3 netRa19 305630.0892935388
Lbr19 netRa19 netL19 1.0364943267394956e-05
Rbbr19 netL19 node_4 1045375.0609088354
Cbr19 netL19 node_4 3.529458174709212e-17

* Branch 20
Rabr20 node_3 netRa20 4493.0137705764455
Lbr20 netRa20 netL20 -4.926528607130883e-07
Rbbr20 netL20 node_4 62508.963214602845
Cbr20 netL20 node_4 -9.139726805805309e-16

* Branch 21
Rabr21 node_3 netRa21 7916902.236617085
Lbr21 netRa21 netL21 2.8455242300608357e-05
Rbbr21 netL21 node_4 8179021.454737164
Cbr21 netL21 node_4 4.444675102580166e-19

* Branch 22
Rabr22 node_3 netRa22 -30923.90600921787
Lbr22 netRa22 netL22 -2.9809810115416195e-07
Rbbr22 netL22 node_4 -39451.700661915325
Cbr22 netL22 node_4 -2.7991215314282387e-16

* Branch 23
Rabr23 node_3 netRa23 -103943.98677464617
Lbr23 netRa23 netL23 1.4777510184841592e-06
Rbbr23 netL23 node_4 -165610.92120369695
Cbr23 netL23 node_4 7.891322187636015e-17

* Branch 24
Rabr24 node_3 netRa24 357879.789971262
Lbr24 netRa24 netL24 -6.156683512578756e-06
Rbbr24 netL24 node_4 681591.0216992487
Cbr24 netL24 node_4 -2.4102052584984645e-17

.ends


* Y'44
.subckt yp44 node_4 node_ref
* Branch 0
Rabr0 node_4 netRa0 -452.1487700651417
Lbr0 netRa0 netL0 -1.4885728677078267e-07
Rbbr0 netL0 node_ref 231.64255043068053
Cbr0 netL0 node_ref -5.262276442702259e-13

* Branch 1
Rabr1 node_4 netRa1 -384.30716748988544
Lbr1 netRa1 netL1 6.963341654817459e-07
Rbbr1 netL1 node_ref -31151.53430446576
Cbr1 netL1 node_ref 3.5950450599452097e-14

* Branch 2
Rabr2 node_4 netRa2 3680.0415576978985
Lbr2 netRa2 netL2 -3.3804679709632905e-06
Rbbr2 netL2 node_ref 108527.48846653324
Cbr2 netL2 node_ref -7.239156140682547e-15

* Branch 3
Rabr3 node_4 netRa3 232.66606248516518
Lbr3 netRa3 netL3 4.174780405864241e-07
Rbbr3 netL3 node_ref -65751.30986626429
Cbr3 netL3 node_ref 6.079481894511066e-14

* Branch 4
Rabr4 node_4 netRa4 -410.5699161517149
Lbr4 netRa4 netL4 3.591212144192571e-07
Rbbr4 netL4 node_ref -4108.259873584922
Cbr4 netL4 node_ref 6.213279729205845e-14

* Branch 5
Rabr5 node_4 netRa5 -1600.178454365244
Lbr5 netRa5 netL5 -1.3635817448866234e-07
Rbbr5 netL5 node_ref -5875.130023194041
Cbr5 netL5 node_ref -4.5663785981364055e-14

* Branch 6
Rabr6 node_4 netRa6 71651.5487257445
Lbr6 netRa6 netL6 -1.4756051698454795e-05
Rbbr6 netL6 node_ref 459449.48027098004
Cbr6 netL6 node_ref -3.6268654899702983e-16

* Branch 7
Rabr7 node_4 netRa7 -296689.5531137229
Lbr7 netRa7 netL7 4.146281646380012e-05
Rbbr7 netL7 node_ref -1151589.179554077
Cbr7 netL7 node_ref 1.1335455222102043e-16

* Branch 8
Rabr8 node_4 netRa8 -91.39343017567465
Lbr8 netRa8 netL8 8.817473395134768e-08
Rbbr8 netL8 node_ref -3301.0010322289554
Cbr8 netL8 node_ref 6.89747807025496e-14

* Branch 9
Rabr9 node_4 netRa9 4482.208444209113
Lbr9 netRa9 netL9 -1.822336140380708e-06
Rbbr9 netL9 node_ref 200406.83802394202
Cbr9 netL9 node_ref -1.5105421899067124e-15

* Branch 10
Rabr10 node_4 netRa10 -32.12322568164358
Lbr10 netRa10 netL10 1.3239485154887825e-07
Rbbr10 netL10 node_ref -31521.41699347519
Cbr10 netL10 node_ref 2.1226807428205986e-14

* Branch 11
Rabr11 node_4 netRa11 13277.961796530944
Lbr11 netRa11 netL11 -4.2641236202950714e-07
Rbbr11 netL11 node_ref 20305.64582304293
Cbr11 netL11 node_ref -1.320007130832125e-15

* Branch 12
Rabr12 node_4 netRa12 606.1244712147017
Lbr12 netRa12 netL12 1.1153893082925438e-07
Rbbr12 netL12 node_ref 16463.673216147286
Cbr12 netL12 node_ref 1.3701002169276064e-14

* Branch 13
Rabr13 node_4 netRa13 -361880.36283068813
Lbr13 netRa13 netL13 -2.334772612953434e-06
Rbbr13 netL13 node_ref -371495.85542881535
Cbr13 netL13 node_ref -1.7547323680098056e-17

* Branch 14
Rabr14 node_4 netRa14 -248.3130592735429
Lbr14 netRa14 netL14 1.0685163613784907e-07
Rbbr14 netL14 node_ref -28615.334500355024
Cbr14 netL14 node_ref 9.388640480927412e-15

* Branch 15
Rabr15 node_4 netRa15 20865.63131764469
Lbr15 netRa15 netL15 7.025772617113829e-07
Rbbr15 netL15 node_ref 46899.280837251536
Cbr15 netL15 node_ref 7.990668977432752e-16

* Branch 16
Rabr16 node_4 netRa16 121.2343241766676
Lbr16 netRa16 netL16 8.540844601562888e-08
Rbbr16 netL16 node_ref -3010019.9823138984
Cbr16 netL16 node_ref 8.24095835418231e-15

* Branch 17
Rabr17 node_4 netRa17 -280415.16917703574
Lbr17 netRa17 netL17 -2.1819550435513953e-06
Rbbr17 netL17 node_ref -305469.3803385434
Cbr17 netL17 node_ref -2.6229943706128355e-17

* Branch 18
Rabr18 node_4 netRa18 37.72490447555568
Lbr18 netRa18 netL18 4.531218463539911e-09
Rbbr18 netL18 node_ref -123.5891455607126
Cbr18 netL18 node_ref 1.8779466995301176e-13

* Branch 19
Rabr19 node_4 netRa19 -13706.713760660063
Lbr19 netRa19 netL19 7.988952679615521e-07
Rbbr19 netL19 node_ref -92789.44149402376
Cbr19 netL19 node_ref 5.515162506461122e-16

* Branch 20
Rabr20 node_4 netRa20 -1334.4181558744956
Lbr20 netRa20 netL20 4.0212975508161237e-08
Rbbr20 netL20 node_ref -3328.514672018788
Cbr20 netL20 node_ref 7.227674818421082e-15

* Branch 21
Rabr21 node_4 netRa21 -539.5122196465381
Lbr21 netRa21 netL21 7.33701760307309e-08
Rbbr21 netL21 node_ref -18251.60225882885
Cbr21 netL21 node_ref 5.2198022013982904e-15

* Branch 22
Rabr22 node_4 netRa22 2109.1353832609666
Lbr22 netRa22 netL22 2.9807929037341016e-08
Rbbr22 netL22 node_ref 3450.3133140889995
Cbr22 netL22 node_ref 5.0339166522824745e-15

* Branch 23
Rabr23 node_4 netRa23 1055.0629981936388
Lbr23 netRa23 netL23 -7.580512212831825e-08
Rbbr23 netL23 node_ref 13099.68720214193
Cbr23 netL23 node_ref -3.798581362513483e-15

* Branch 24
Rabr24 node_4 netRa24 -8865.459020453683
Lbr24 netRa24 netL24 -5.217440564948421e-07
Rbbr24 netL24 node_ref -126067.91774582065
Cbr24 netL24 node_ref -5.567261023845991e-16

.ends


.end
